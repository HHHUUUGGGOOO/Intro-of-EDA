//
// Conformal-LEC Version 19.20-d218 (25-Feb-2020)
//
module top(\A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,
        \A[2][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,
        \A[1][0] ,\A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,
        \A[0][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,
        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ,\O[19] ,
        \O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,\O[10] ,\O[9] ,
        \O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,\O[0] );
input \A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,
        \A[2][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,
        \A[1][0] ,\A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,
        \A[0][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,
        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ;
output \O[19] ,\O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,
        \O[10] ,\O[9] ,\O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,
        \O[0] ;

wire \69_ZERO , \70_ZERO , \71_ZERO , \72_ZERO , \73_ZERO , \74_ZERO , \75_ZERO , \76 , \77 ,
         \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86_ONE , \87_ONE ,
         \88 , \89 , \90 , \91 , \92 , \93 , \94 , \95 , \96 , \97 ,
         \98 , \99 , \100 , \101 , \102 , \103 , \104 , \105 , \106 , \107 ,
         \108 , \109_A[9] , \110 , \111 , \112 , \113 , \114 , \115_A[8] , \116 , \117 ,
         \118 , \119 , \120 , \121_A[7] , \122 , \123 , \124 , \125 , \126 , \127_A[6] ,
         \128 , \129 , \130 , \131 , \132 , \133_A[5] , \134 , \135 , \136 , \137 ,
         \138 , \139_A[4] , \140 , \141 , \142 , \143 , \144 , \145_A[3] , \146 , \147 ,
         \148 , \149 , \150 , \151_A[2] , \152 , \153 , \154 , \155 , \156 , \157_A[1] ,
         \158 , \159 , \160 , \161 , \162 , \163_A[0] , \164_B[9] , \165_B[8] , \166_B[7] , \167_B[6] ,
         \168_B[5] , \169_B[4] , \170_B[3] , \171_B[2] , \172_B[1] , \173_B[0] , \174 , \175 , \176 , \177 ,
         \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 ,
         \188 , \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 ,
         \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 ,
         \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 ,
         \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 ,
         \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 ,
         \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 ,
         \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 ,
         \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 ,
         \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 ,
         \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 ,
         \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 ,
         \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 ,
         \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 ,
         \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 ,
         \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 ,
         \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 ,
         \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 ,
         \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 ,
         \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 ,
         \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 ,
         \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 ,
         \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 ,
         \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 ,
         \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 ,
         \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 ,
         \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 ,
         \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 ,
         \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 ,
         \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 ,
         \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 ,
         \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 ,
         \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 ,
         \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 ,
         \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 ,
         \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 ,
         \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 ,
         \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 ,
         \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 ,
         \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 ,
         \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 ,
         \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 ,
         \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 ,
         \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 ,
         \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 ,
         \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 ,
         \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 ,
         \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,
         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,
         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675_Z[19] , \676 , \677_Z[18] ,
         \678 , \679_Z[17] , \680 , \681_Z[16] , \682 , \683_Z[15] , \684 , \685_Z[14] , \686 , \687_Z[13] ,
         \688 , \689_Z[12] , \690 , \691_Z[11] , \692 , \693_Z[10] , \694 , \695_Z[9] , \696 , \697_Z[8] ,
         \698 , \699_Z[7] , \700 , \701_Z[6] , \702 , \703_Z[5] , \704 , \705_Z[4] , \706 , \707_Z[3] ,
         \708 , \709_Z[2] , \710 , \711_Z[1] , \712 , \713_Z[0] ;
buf ( \O[19] , \675_Z[19] );
buf ( \O[18] , \677_Z[18] );
buf ( \O[17] , \679_Z[17] );
buf ( \O[16] , \681_Z[16] );
buf ( \O[15] , \683_Z[15] );
buf ( \O[14] , \685_Z[14] );
buf ( \O[13] , \687_Z[13] );
buf ( \O[12] , \689_Z[12] );
buf ( \O[11] , \691_Z[11] );
buf ( \O[10] , \693_Z[10] );
buf ( \O[9] , \695_Z[9] );
buf ( \O[8] , \697_Z[8] );
buf ( \O[7] , \699_Z[7] );
buf ( \O[6] , \701_Z[6] );
buf ( \O[5] , \703_Z[5] );
buf ( \O[4] , \705_Z[4] );
buf ( \O[3] , \707_Z[3] );
buf ( \O[2] , \709_Z[2] );
buf ( \O[1] , \711_Z[1] );
buf ( \O[0] , \713_Z[0] );
not ( \88 , \I[1] );
nor ( \89 , \I[0] , \88 , \I[2] , \I[3] , \I[4] , \I[5] , \I[6] , \I[7] );
and ( \90 , \A[2][9] , \89 );
not ( \91 , \I[0] );
nor ( \92 , \91 , \I[1] , \I[2] , \I[3] , \I[4] , \I[5] , \I[6] , \I[7] );
and ( \93 , \A[1][9] , \92 );
nor ( \94 , \I[0] , \I[1] , \I[2] , \I[3] , \I[4] , \I[5] , \I[6] , \I[7] );
and ( \95 , \A[0][9] , \94 );
or ( \96 , \90 , \93 , \95 );
buf ( \97 , \I[2] );
buf ( \98 , \I[3] );
buf ( \99 , \I[4] );
buf ( \100 , \I[5] );
buf ( \101 , \I[6] );
buf ( \102 , \I[7] );
buf ( \103 , \I[1] );
buf ( \104 , \I[0] );
and ( \105 , \103 , \104 );
or ( \106 , \97 , \98 , \99 , \100 , \101 , \102 , \105 );
buf ( \107 , \106 );
_DC ( \108 , \96 , \107 );
buf ( \109_A[9] , \108 );
and ( \110 , \A[2][8] , \89 );
and ( \111 , \A[1][8] , \92 );
and ( \112 , \A[0][8] , \94 );
or ( \113 , \110 , \111 , \112 );
_DC ( \114 , \113 , \107 );
buf ( \115_A[8] , \114 );
and ( \116 , \A[2][7] , \89 );
and ( \117 , \A[1][7] , \92 );
and ( \118 , \A[0][7] , \94 );
or ( \119 , \116 , \117 , \118 );
_DC( \120 , \119 , \107 );
buf ( \121_A[7] , \120 );
and ( \122 , \A[2][6] , \89 );
and ( \123 , \A[1][6] , \92 );
and ( \124 , \A[0][6] , \94 );
or ( \125 , \122 , \123 , \124 );
_DC ( \126 , \125 , \107 );
buf ( \127_A[6] , \126 );
and ( \128 , \A[2][5] , \89 );
and ( \129 , \A[1][5] , \92 );
and ( \130 , \A[0][5] , \94 );
or ( \131 , \128 , \129 , \130 );
_DC ( \132 , \131 , \107 );
buf ( \133_A[5] , \132 );
and ( \134 , \A[2][4] , \89 );
and ( \135 , \A[1][4] , \92 );
and ( \136 , \A[0][4] , \94 );
or ( \137 , \134 , \135 , \136 );
_DC ( \138 , \137 , \107 );
buf ( \139_A[4] , \138 );
and ( \140 , \A[2][3] , \89 );
and ( \141 , \A[1][3] , \92 );
and ( \142 , \A[0][3] , \94 );
or ( \143 , \140 , \141 , \142 );
_DC ( \144 , \143 , \107 );
buf ( \145_A[3] , \144 );
and ( \146 , \A[2][2] , \89 );
and ( \147 , \A[1][2] , \92 );
and ( \148 , \A[0][2] , \94 );
or ( \149 , \146 , \147 , \148 );
_DC ( \150 , \149 , \107 );
buf ( \151_A[2] , \150 );
and ( \152 , \A[2][1] , \89 );
and ( \153 , \A[1][1] , \92 );
and ( \154 , \A[0][1] , \94 );
or ( \155 , \152 , \153 , \154 );
_DC ( \156 , \155 , \107 );
buf ( \157_A[1] , \156 );
and ( \158 , \A[2][0] , \89 );
and ( \159 , \A[1][0] , \92 );
and ( \160 , \A[0][0] , \94 );
or ( \161 , \158 , \159 , \160 );
_DC ( \162 , \161 , \107 );
buf ( \163_A[0] , \162 );
buf ( \164_B[9] , \B[9] );
buf ( \165_B[8] , \B[8] );
buf ( \166_B[7] , \B[7] );
buf ( \167_B[6] , \B[6] );
buf ( \168_B[5] , \B[5] );
buf ( \169_B[4] , \B[4] );
buf ( \170_B[3] , \B[3] );
buf ( \171_B[2] , \B[2] );
buf ( \172_B[1] , \B[1] );
buf ( \173_B[0] , \B[0] );
and ( \174 , \109_A[9] , \172_B[1] );
and ( \175 , \109_A[9] , \173_B[0] );
and ( \176 , \115_A[8] , \172_B[1] );
and ( \177 , \175 , \176 );
xor ( \178 , \175 , \176 );
and ( \179 , \115_A[8] , \173_B[0] );
and ( \180 , \121_A[7] , \172_B[1] );
and ( \181 , \179 , \180 );
xor ( \182 , \179 , \180 );
and ( \183 , \121_A[7] , \173_B[0] );
and ( \184 , \127_A[6] , \172_B[1] );
and ( \185 , \183 , \184 );
xor ( \186 , \183 , \184 );
and ( \187 , \127_A[6] , \173_B[0] );
and ( \188 , \133_A[5] , \172_B[1] );
and ( \189 , \187 , \188 );
xor ( \190 , \187 , \188 );
and ( \191 , \133_A[5] , \173_B[0] );
and ( \192 , \139_A[4] , \172_B[1] );
and ( \193 , \191 , \192 );
xor ( \194 , \191 , \192 );
and ( \195 , \139_A[4] , \173_B[0] );
and ( \196 , \145_A[3] , \172_B[1] );
and ( \197 , \195 , \196 );
xor ( \198 , \195 , \196 );
and ( \199 , \145_A[3] , \173_B[0] );
and ( \200 , \151_A[2] , \172_B[1] );
and ( \201 , \199 , \200 );
xor ( \202 , \199 , \200 );
and ( \203 , \151_A[2] , \173_B[0] );
and ( \204 , \157_A[1] , \172_B[1] );
and ( \205 , \203 , \204 );
xor ( \206 , \203 , \204 );
and ( \207 , \157_A[1] , \173_B[0] );
and ( \208 , \163_A[0] , \172_B[1] );
and ( \209 , \207 , \208 );
and ( \210 , \206 , \209 );
or ( \211 , \205 , \210 );
and ( \212 , \202 , \211 );
or ( \213 , \201 , \212 );
and ( \214 , \198 , \213 );
or ( \215 , \197 , \214 );
and ( \216 , \194 , \215 );
or ( \217 , \193 , \216 );
and ( \218 , \190 , \217 );
or ( \219 , \189 , \218 );
and ( \220 , \186 , \219 );
or ( \221 , \185 , \220 );
and ( \222 , \182 , \221 );
or ( \223 , \181 , \222 );
and ( \224 , \178 , \223 );
or ( \225 , \177 , \224 );
and ( \226 , \174 , \225 );
and ( \227 , \109_A[9] , \171_B[2] );
and ( \228 , \226 , \227 );
xor ( \229 , \226 , \227 );
xor ( \230 , \174 , \225 );
and ( \231 , \115_A[8] , \171_B[2] );
and ( \232 , \230 , \231 );
xor ( \233 , \230 , \231 );
xor ( \234 , \178 , \223 );
and ( \235 , \121_A[7] , \171_B[2] );
and ( \236 , \234 , \235 );
xor ( \237 , \234 , \235 );
xor ( \238 , \182 , \221 );
and ( \239 , \127_A[6] , \171_B[2] );
and ( \240 , \238 , \239 );
xor ( \241 , \238 , \239 );
xor ( \242 , \186 , \219 );
and ( \243 , \133_A[5] , \171_B[2] );
and ( \244 , \242 , \243 );
xor ( \245 , \242 , \243 );
xor ( \246 , \190 , \217 );
and ( \247 , \139_A[4] , \171_B[2] );
and ( \248 , \246 , \247 );
xor ( \249 , \246 , \247 );
xor ( \250 , \194 , \215 );
and ( \251 , \145_A[3] , \171_B[2] );
and ( \252 , \250 , \251 );
xor ( \253 , \250 , \251 );
xor ( \254 , \198 , \213 );
and ( \255 , \151_A[2] , \171_B[2] );
and ( \256 , \254 , \255 );
xor ( \257 , \254 , \255 );
xor ( \258 , \202 , \211 );
and ( \259 , \157_A[1] , \171_B[2] );
and ( \260 , \258 , \259 );
xor ( \261 , \258 , \259 );
xor ( \262 , \206 , \209 );
and ( \263 , \163_A[0] , \171_B[2] );
and ( \264 , \262 , \263 );
and ( \265 , \261 , \264 );
or ( \266 , \260 , \265 );
and ( \267 , \257 , \266 );
or ( \268 , \256 , \267 );
and ( \269 , \253 , \268 );
or ( \270 , \252 , \269 );
and ( \271 , \249 , \270 );
or ( \272 , \248 , \271 );
and ( \273 , \245 , \272 );
or ( \274 , \244 , \273 );
and ( \275 , \241 , \274 );
or ( \276 , \240 , \275 );
and ( \277 , \237 , \276 );
or ( \278 , \236 , \277 );
and ( \279 , \233 , \278 );
or ( \280 , \232 , \279 );
and ( \281 , \229 , \280 );
or ( \282 , \228 , \281 );
and ( \283 , \109_A[9] , \170_B[3] );
and ( \284 , \282 , \283 );
xor ( \285 , \282 , \283 );
xor ( \286 , \229 , \280 );
and ( \287 , \115_A[8] , \170_B[3] );
and ( \288 , \286 , \287 );
xor ( \289 , \286 , \287 );
xor ( \290 , \233 , \278 );
and ( \291 , \121_A[7] , \170_B[3] );
and ( \292 , \290 , \291 );
xor ( \293 , \290 , \291 );
xor ( \294 , \237 , \276 );
and ( \295 , \127_A[6] , \170_B[3] );
and ( \296 , \294 , \295 );
xor ( \297 , \294 , \295 );
xor ( \298 , \241 , \274 );
and ( \299 , \133_A[5] , \170_B[3] );
and ( \300 , \298 , \299 );
xor ( \301 , \298 , \299 );
xor ( \302 , \245 , \272 );
and ( \303 , \139_A[4] , \170_B[3] );
and ( \304 , \302 , \303 );
xor ( \305 , \302 , \303 );
xor ( \306 , \249 , \270 );
and ( \307 , \145_A[3] , \170_B[3] );
and ( \308 , \306 , \307 );
xor ( \309 , \306 , \307 );
xor ( \310 , \253 , \268 );
and ( \311 , \151_A[2] , \170_B[3] );
and ( \312 , \310 , \311 );
xor ( \313 , \310 , \311 );
xor ( \314 , \257 , \266 );
and ( \315 , \157_A[1] , \170_B[3] );
and ( \316 , \314 , \315 );
xor ( \317 , \314 , \315 );
xor ( \318 , \261 , \264 );
and ( \319 , \163_A[0] , \170_B[3] );
and ( \320 , \318 , \319 );
and ( \321 , \317 , \320 );
or ( \322 , \316 , \321 );
and ( \323 , \313 , \322 );
or ( \324 , \312 , \323 );
and ( \325 , \309 , \324 );
or ( \326 , \308 , \325 );
and ( \327 , \305 , \326 );
or ( \328 , \304 , \327 );
and ( \329 , \301 , \328 );
or ( \330 , \300 , \329 );
and ( \331 , \297 , \330 );
or ( \332 , \296 , \331 );
and ( \333 , \293 , \332 );
or ( \334 , \292 , \333 );
and ( \335 , \289 , \334 );
or ( \336 , \288 , \335 );
and ( \337 , \285 , \336 );
or ( \338 , \284 , \337 );
and ( \339 , \109_A[9] , \169_B[4] );
and ( \340 , \338 , \339 );
xor ( \341 , \338 , \339 );
xor ( \342 , \285 , \336 );
and ( \343 , \115_A[8] , \169_B[4] );
and ( \344 , \342 , \343 );
xor ( \345 , \342 , \343 );
xor ( \346 , \289 , \334 );
and ( \347 , \121_A[7] , \169_B[4] );
and ( \348 , \346 , \347 );
xor ( \349 , \346 , \347 );
xor ( \350 , \293 , \332 );
and ( \351 , \127_A[6] , \169_B[4] );
and ( \352 , \350 , \351 );
xor ( \353 , \350 , \351 );
xor ( \354 , \297 , \330 );
and ( \355 , \133_A[5] , \169_B[4] );
and ( \356 , \354 , \355 );
xor ( \357 , \354 , \355 );
xor ( \358 , \301 , \328 );
and ( \359 , \139_A[4] , \169_B[4] );
and ( \360 , \358 , \359 );
xor ( \361 , \358 , \359 );
xor ( \362 , \305 , \326 );
and ( \363 , \145_A[3] , \169_B[4] );
and ( \364 , \362 , \363 );
xor ( \365 , \362 , \363 );
xor ( \366 , \309 , \324 );
and ( \367 , \151_A[2] , \169_B[4] );
and ( \368 , \366 , \367 );
xor ( \369 , \366 , \367 );
xor ( \370 , \313 , \322 );
and ( \371 , \157_A[1] , \169_B[4] );
and ( \372 , \370 , \371 );
xor ( \373 , \370 , \371 );
xor ( \374 , \317 , \320 );
and ( \375 , \163_A[0] , \169_B[4] );
and ( \376 , \374 , \375 );
and ( \377 , \373 , \376 );
or ( \378 , \372 , \377 );
and ( \379 , \369 , \378 );
or ( \380 , \368 , \379 );
and ( \381 , \365 , \380 );
or ( \382 , \364 , \381 );
and ( \383 , \361 , \382 );
or ( \384 , \360 , \383 );
and ( \385 , \357 , \384 );
or ( \386 , \356 , \385 );
and ( \387 , \353 , \386 );
or ( \388 , \352 , \387 );
and ( \389 , \349 , \388 );
or ( \390 , \348 , \389 );
and ( \391 , \345 , \390 );
or ( \392 , \344 , \391 );
and ( \393 , \341 , \392 );
or ( \394 , \340 , \393 );
and ( \395 , \109_A[9] , \168_B[5] );
and ( \396 , \394 , \395 );
xor ( \397 , \394 , \395 );
xor ( \398 , \341 , \392 );
and ( \399 , \115_A[8] , \168_B[5] );
and ( \400 , \398 , \399 );
xor ( \401 , \398 , \399 );
xor ( \402 , \345 , \390 );
and ( \403 , \121_A[7] , \168_B[5] );
and ( \404 , \402 , \403 );
xor ( \405 , \402 , \403 );
xor ( \406 , \349 , \388 );
and ( \407 , \127_A[6] , \168_B[5] );
and ( \408 , \406 , \407 );
xor ( \409 , \406 , \407 );
xor ( \410 , \353 , \386 );
and ( \411 , \133_A[5] , \168_B[5] );
and ( \412 , \410 , \411 );
xor ( \413 , \410 , \411 );
xor ( \414 , \357 , \384 );
and ( \415 , \139_A[4] , \168_B[5] );
and ( \416 , \414 , \415 );
xor ( \417 , \414 , \415 );
xor ( \418 , \361 , \382 );
and ( \419 , \145_A[3] , \168_B[5] );
and ( \420 , \418 , \419 );
xor ( \421 , \418 , \419 );
xor ( \422 , \365 , \380 );
and ( \423 , \151_A[2] , \168_B[5] );
and ( \424 , \422 , \423 );
xor ( \425 , \422 , \423 );
xor ( \426 , \369 , \378 );
and ( \427 , \157_A[1] , \168_B[5] );
and ( \428 , \426 , \427 );
xor ( \429 , \426 , \427 );
xor ( \430 , \373 , \376 );
and ( \431 , \163_A[0] , \168_B[5] );
and ( \432 , \430 , \431 );
and ( \433 , \429 , \432 );
or ( \434 , \428 , \433 );
and ( \435 , \425 , \434 );
or ( \436 , \424 , \435 );
and ( \437 , \421 , \436 );
or ( \438 , \420 , \437 );
and ( \439 , \417 , \438 );
or ( \440 , \416 , \439 );
and ( \441 , \413 , \440 );
or ( \442 , \412 , \441 );
and ( \443 , \409 , \442 );
or ( \444 , \408 , \443 );
and ( \445 , \405 , \444 );
or ( \446 , \404 , \445 );
and ( \447 , \401 , \446 );
or ( \448 , \400 , \447 );
and ( \449 , \397 , \448 );
or ( \450 , \396 , \449 );
and ( \451 , \109_A[9] , \167_B[6] );
and ( \452 , \450 , \451 );
xor ( \453 , \450 , \451 );
xor ( \454 , \397 , \448 );
and ( \455 , \115_A[8] , \167_B[6] );
and ( \456 , \454 , \455 );
xor ( \457 , \454 , \455 );
xor ( \458 , \401 , \446 );
and ( \459 , \121_A[7] , \167_B[6] );
and ( \460 , \458 , \459 );
xor ( \461 , \458 , \459 );
xor ( \462 , \405 , \444 );
and ( \463 , \127_A[6] , \167_B[6] );
and ( \464 , \462 , \463 );
xor ( \465 , \462 , \463 );
xor ( \466 , \409 , \442 );
and ( \467 , \133_A[5] , \167_B[6] );
and ( \468 , \466 , \467 );
xor ( \469 , \466 , \467 );
xor ( \470 , \413 , \440 );
and ( \471 , \139_A[4] , \167_B[6] );
and ( \472 , \470 , \471 );
xor ( \473 , \470 , \471 );
xor ( \474 , \417 , \438 );
and ( \475 , \145_A[3] , \167_B[6] );
and ( \476 , \474 , \475 );
xor ( \477 , \474 , \475 );
xor ( \478 , \421 , \436 );
and ( \479 , \151_A[2] , \167_B[6] );
and ( \480 , \478 , \479 );
xor ( \481 , \478 , \479 );
xor ( \482 , \425 , \434 );
and ( \483 , \157_A[1] , \167_B[6] );
and ( \484 , \482 , \483 );
xor ( \485 , \482 , \483 );
xor ( \486 , \429 , \432 );
and ( \487 , \163_A[0] , \167_B[6] );
and ( \488 , \486 , \487 );
and ( \489 , \485 , \488 );
or ( \490 , \484 , \489 );
and ( \491 , \481 , \490 );
or ( \492 , \480 , \491 );
and ( \493 , \477 , \492 );
or ( \494 , \476 , \493 );
and ( \495 , \473 , \494 );
or ( \496 , \472 , \495 );
and ( \497 , \469 , \496 );
or ( \498 , \468 , \497 );
and ( \499 , \465 , \498 );
or ( \500 , \464 , \499 );
and ( \501 , \461 , \500 );
or ( \502 , \460 , \501 );
and ( \503 , \457 , \502 );
or ( \504 , \456 , \503 );
and ( \505 , \453 , \504 );
or ( \506 , \452 , \505 );
and ( \507 , \109_A[9] , \166_B[7] );
and ( \508 , \506 , \507 );
xor ( \509 , \506 , \507 );
xor ( \510 , \453 , \504 );
and ( \511 , \115_A[8] , \166_B[7] );
and ( \512 , \510 , \511 );
xor ( \513 , \510 , \511 );
xor ( \514 , \457 , \502 );
and ( \515 , \121_A[7] , \166_B[7] );
and ( \516 , \514 , \515 );
xor ( \517 , \514 , \515 );
xor ( \518 , \461 , \500 );
and ( \519 , \127_A[6] , \166_B[7] );
and ( \520 , \518 , \519 );
xor ( \521 , \518 , \519 );
xor ( \522 , \465 , \498 );
and ( \523 , \133_A[5] , \166_B[7] );
and ( \524 , \522 , \523 );
xor ( \525 , \522 , \523 );
xor ( \526 , \469 , \496 );
and ( \527 , \139_A[4] , \166_B[7] );
and ( \528 , \526 , \527 );
xor ( \529 , \526 , \527 );
xor ( \530 , \473 , \494 );
and ( \531 , \145_A[3] , \166_B[7] );
and ( \532 , \530 , \531 );
xor ( \533 , \530 , \531 );
xor ( \534 , \477 , \492 );
and ( \535 , \151_A[2] , \166_B[7] );
and ( \536 , \534 , \535 );
xor ( \537 , \534 , \535 );
xor ( \538 , \481 , \490 );
and ( \539 , \157_A[1] , \166_B[7] );
and ( \540 , \538 , \539 );
xor ( \541 , \538 , \539 );
xor ( \542 , \485 , \488 );
and ( \543 , \163_A[0] , \166_B[7] );
and ( \544 , \542 , \543 );
and ( \545 , \541 , \544 );
or ( \546 , \540 , \545 );
and ( \547 , \537 , \546 );
or ( \548 , \536 , \547 );
and ( \549 , \533 , \548 );
or ( \550 , \532 , \549 );
and  ( \551 , \529 , \550 );
or  ( \552 , \528 , \551 );
and  ( \553 , \525 , \552 );
or  ( \554 , \524 , \553 );
and ( \555 , \521 , \554 );
or ( \556 , \520 , \555 );
and  ( \557 , \517 , \556 );
or  ( \558 , \516 , \557 );
and  ( \559 , \513 , \558 );
or  ( \560 , \512 , \559 );
and  ( \561 , \509 , \560 );
or  ( \562 , \508 , \561 );
and  ( \563 , \109_A[9] , \165_B[8] );
and ( \564 , \562 , \563 );
xor ( \565 , \562 , \563 );
xor ( \566 , \509 , \560 );
and  ( \567 , \115_A[8] , \165_B[8] );
and ( \568 , \566 , \567 );
xor ( \569 , \566 , \567 );
xor ( \570 , \513 , \558 );
and ( \571 , \121_A[7] , \165_B[8] );
and ( \572 , \570 , \571 );
xor ( \573 , \570 , \571 );
xor ( \574 , \517 , \556 );
and ( \575 , \127_A[6] , \165_B[8] );
and ( \576 , \574 , \575 );
xor ( \577 , \574 , \575 );
xor ( \578 , \521 , \554 );
and ( \579 , \133_A[5] , \165_B[8] );
and ( \580 , \578 , \579 );
xor ( \581 , \578 , \579 );
xor ( \582 , \525 , \552 );
and ( \583 , \139_A[4] , \165_B[8] );
and ( \584 , \582 , \583 );
xor ( \585 , \582 , \583 );
xor ( \586 , \529 , \550 );
and ( \587 , \145_A[3] , \165_B[8] );
and ( \588 , \586 , \587 );
xor ( \589 , \586 , \587 );
xor ( \590 , \533 , \548 );
and ( \591 , \151_A[2] , \165_B[8] );
and ( \592 , \590 , \591 );
xor ( \593 , \590 , \591 );
xor ( \594 , \537 , \546 );
and ( \595 , \157_A[1] , \165_B[8] );
and ( \596 , \594 , \595 );
xor ( \597 , \594 , \595 );
xor ( \598 , \541 , \544 );
and ( \599 , \163_A[0] , \165_B[8] );
and ( \600 , \598 , \599 );
and ( \601 , \597 , \600 );
or  ( \602 , \596 , \601 );
and ( \603 , \593 , \602 );
or ( \604 , \592 , \603 );
and ( \605 , \589 , \604 );
or ( \606 , \588 , \605 );
and ( \607 , \585 , \606 );
or ( \608 , \584 , \607 );
and ( \609 , \581 , \608 );
or ( \610 , \580 , \609 );
and ( \611 , \577 , \610 );
or ( \612 , \576 , \611 );
and ( \613 , \573 , \612 );
or ( \614 , \572 , \613 );
and ( \615 , \569 , \614 );
or ( \616 , \568 , \615 );
and ( \617 , \565 , \616 );
or ( \618 , \564 , \617 );
and ( \619 , \109_A[9] , \164_B[9] );
and ( \620 , \618 , \619 );
xor ( \621 , \618 , \619 );
xor ( \622 , \565 , \616 );
and ( \623 , \115_A[8] , \164_B[9] );
and ( \624 , \622 , \623 );
xor ( \625 , \622 , \623 );
xor ( \626 , \569 , \614 );
and ( \627 , \121_A[7] , \164_B[9] );
and ( \628 , \626 , \627 );
xor ( \629 , \626 , \627 );
xor ( \630 , \573 , \612 );
and ( \631 , \127_A[6] , \164_B[9] );
and ( \632 , \630 , \631 );
xor ( \633 , \630 , \631 );
xor ( \634 , \577 , \610 );
and ( \635 , \133_A[5] , \164_B[9] );
and ( \636 , \634 , \635 );
xor ( \637 , \634 , \635 );
xor ( \638 , \581 , \608 );
and ( \639 , \139_A[4] , \164_B[9] );
and ( \640 , \638 , \639 );
xor ( \641 , \638 , \639 );
xor ( \642 , \585 , \606 );
and ( \643 , \145_A[3] , \164_B[9] );
and ( \644 , \642 , \643 );
xor ( \645 , \642 , \643 );
xor ( \646 , \589 , \604 );
and ( \647 , \151_A[2] , \164_B[9] );
and ( \648 , \646 , \647 );
xor ( \649 , \646 , \647 );
xor ( \650 , \593 , \602 );
and ( \651 , \157_A[1] , \164_B[9] );
and ( \652 , \650 , \651 );
xor ( \653 , \650 , \651 );
xor ( \654 , \597 , \600 );
and ( \655 , \163_A[0] , \164_B[9] );
and ( \656 , \654 , \655 );
and ( \657 , \653 , \656 );
or ( \658 , \652 , \657 );
and ( \659 , \649 , \658 );
or ( \660 , \648 , \659 );
and ( \661 , \645 , \660 );
or ( \662 , \644 , \661 );
and ( \663 , \641 , \662 );
or ( \664 , \640 , \663 );
and ( \665 , \637 , \664 );
or ( \666 , \636 , \665 );
and ( \667 , \633 , \666 );
or ( \668 , \632 , \667 );
and ( \669 , \629 , \668 );
or ( \670 , \628 , \669 );
and ( \671 , \625 , \670 );
or ( \672 , \624 , \671 );
and ( \673 , \621 , \672 );
or ( \674 , \620 , \673 );
buf ( \675_Z[19] , \674 );
xor ( \676 , \621 , \672 );
buf ( \677_Z[18] , \676 );
xor ( \678 , \625 , \670 );
buf ( \679_Z[17] , \678 );
xor ( \680 , \629 , \668 );
buf ( \681_Z[16] , \680 );
xor ( \682 , \633 , \666 );
buf ( \683_Z[15] , \682 );
xor ( \684 , \637 , \664 );
buf ( \685_Z[14] , \684 );
xor ( \686 , \641 , \662 );
buf ( \687_Z[13] , \686 );
xor ( \688 , \645 , \660 );
buf ( \689_Z[12] , \688 );
xor ( \690 , \649 , \658 );
buf ( \691_Z[11] , \690 );
xor ( \692 , \653 , \656 );
buf ( \693_Z[10] , \692 );
xor ( \694 , \654 , \655 );
buf ( \695_Z[9] , \694 );
xor ( \696 , \598 , \599 );
buf ( \697_Z[8] , \696 );
xor ( \698 , \542 , \543 );
buf ( \699_Z[7] , \698 );
xor ( \700 , \486 , \487 );
buf ( \701_Z[6] , \700 );
xor ( \702 , \430 , \431 );
buf ( \703_Z[5] , \702 );
xor ( \704 , \374 , \375 );
buf ( \705_Z[4] , \704 );
xor ( \706 , \318 , \319 );
buf ( \707_Z[3] , \706 );
xor ( \708 , \262 , \263 );
buf ( \709_Z[2] , \708 );
xor ( \710 , \207 , \208 );
buf ( \711_Z[1] , \710 );
and ( \712 , \163_A[0] , \173_B[0] );
buf ( \713_Z[0] , \712 );
endmodule
